-- MIT License
--
-- Copyright (c) 2019 Oliver Knodel
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE. 

--
-- Author: Oliver Knodel <oliver.knodel@mailbox.tu-dresden.de>
-- Project:	FPGA-DNA-Sequence-Search
--
-- Gather tree with an or in every bode.
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity gather_or_tree is
	generic(
		MODULES			: positive := 512
	);
   Port ( 
		clk 					: in  STD_LOGIC;
		gather_data_in 	: in  STD_LOGIC_VECTOR((MODULES-1) downto 0);
      gather_data_out	: out STD_LOGIC
	);
end gather_or_tree;

architecture Behavioral of gather_or_tree is

	function min(arg1 : integer; arg2 : integer) return integer is
	begin
		if arg1 < arg2 then 
			return arg1; 
		else
			return arg2;
		end if;
	end;

	function node2level(arg : positive) return natural is
		variable tmp : positive;
		variable log : natural;
	begin
		if arg = 1 then
			return 1;
		end if;
    
		tmp := 1;
		log := 1;

		while arg > tmp-1 loop
			tmp := tmp * 2;
			log := log + 1;
		end loop;
		return log-1;
	end;

begin

	gather: block

		constant D 			: positive := 2;-- Node Fan in/out must be 2!
		constant M 			: positive := 1+((MODULES-2)/(D-1)); --internal node count

		signal tree			: std_logic_vector(0 to (M+MODULES-1));
		
			
	begin
		--root connection
		gather_data_out <= tree(0);

		--generate leaves 
		genLeaves: for b in 0 to MODULES-1 generate
			tree(M+b) 		<= gather_data_in(b);
		end generate genLeaves;

		--internal nodes
		genNodes: for b in 0 to M-1 generate
			constant CHILD_FIRST : positive 	:= D*b+1;
			constant CHILD_LAST 	: positive 	:= min(D*b+D, M+MODULES-1);
			constant LEVEL 		: integer 	:= node2level(b+1)-1;
				
			signal node_in_1	: std_logic;
			signal node_in_2	: std_logic;
			signal node_out	: std_logic;

			
		begin
		
			node_in_1 	<= tree(CHILD_FIRST);
			node_in_2 	<= tree(CHILD_LAST);
			
			node_out <= node_in_1 or node_in_2;
			
				process(clk)
				begin
					if rising_edge(clk) then
						tree(b) 		 <= node_out;
					end if;
				end process;
 

		end generate genNodes;
		
	end block gather;

end Behavioral;
